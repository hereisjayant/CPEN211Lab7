
//NOTE: Instance name of your memory is MEM for the auto-grader.


module lab7_top(KEY,SW,LEDR,HEX0,HEX1,HEX2,HEX3,HEX4,HEX5);
  input [3:0] KEY;
  input [9:0] SW;
  output [9:0] LEDR;
  output [6:0] HEX0, HEX1, HEX2, HEX3, HEX4, HEX5;

//------------------------------------------------------------------------------

//Wires:


//------------------------------------------------------------------------------

//Declared modules:

  cpu CPU(clk, reset, read_data, mem_cmd, mem_addr, out, N, V, Z);
  
